/**********************************************************************
 *
 * Vector Space System Project / Material Library Module / IAPWS-IF97
 *
 * Copyright (C) 2020 CIAE.
 *
 * This is free software; you can redistribute and/or modify it under
 * the terms of the GNU Lesser General Public Licence as published
 * by the Free Software Foundation.
 * See the COPYING file for more information.
 *
 * File: common.v
 * Author: YU YANG
 * Created Time: 2020-05-07
 * Version: 0.0.1
 *
 **********************************************************************/
module if97

//****************************************************************
/* Constants used throughout IAPWS-IF97 */
//****************************************************************
const (
	if97_pmax = 100.0  		/* MPa */
	if97_tmin = 273.15 		/* K */
	if97_tmax = 1073.15 		/* K */
	if97_tcrit = 647.096 	/* K */
	if97_pcrit = 22.064 		/* MPa */
	if97_rhocrit = 322.0		/* kg/m³ */
	if97_ptriple = 611.657 	/* Pa */
	if97_r = 0.461526 		/* kJ/kgK */
)

const (
	// Region1
	tmax_region1 = 623.15 		/* K */
	pstar_region1 = 16.53	 	/* MPa */
	tstar_region1 = 1386.0 		/* K */
	// Region2
	tmax_region2 = 1073.15 		/* K */
	tstar_region2 = 540.0 		/* K */
	// Region3
	rhostar_region3 = 322.0		/* kg/m3 */
	tstar_region3 = 647.096		/* K */
	// Region4
	tstar_region4 = 1.0 			/* K */
	// Region5
	tstar_region5 = 1000.0 		/* K */
	// Common
	pstar_region245 = 1.0	 	/* MPa */
)

/* Data struct used throughout IAPWS-IF97 */
struct IJN{
	i_ int
	j_ int
	n_ f64
}

struct FIJN{
	i_ f64
	j_ int
	n_ f64
}

struct JN{
	j_ int
	n_ f64
}

fn ijn(i int,j int,n f64) IJN {	return IJN{i_:i, j_:j, n_:n} }
fn fijn(i f64,j int,n f64) FIJN { return FIJN{i_:i, j_:j, n_:n} }
fn jn(j int,n f64) JN { return JN{j_:j, n_:n} }


//****************************************************************
// CONST FOR `REGION` EQUATIONS
//****************************************************************
const(
	// Region1
	pt_r1 = [	ijn(0, -2, 0.14632971213167E+00),
				ijn(0, -1, -0.84548187169114E+00),
				ijn(0, 0, -0.37563603672040E+01),
				ijn(0, 1, 0.33855169168385E+01),
				ijn(0, 2, -0.95791963387872E+00),
				ijn(0, 3, 0.15772038513228E+00),
				ijn(0, 4, -0.16616417199501E-01),
				ijn(0, 5, 0.81214629983568E-03),
				ijn(1, -9, 0.28319080123804E-03),
				ijn(1, -7, -0.60706301565874E-03),
				ijn(1, -1, -0.18990068218419E-01),
				ijn(1, 0, -0.32529748770505E-01),
				ijn(1, 1, -0.21841717175414E-01),
				ijn(1, 3, -0.52838357969930E-04),
				ijn(2, -3, -0.47184321073267E-03),
				ijn(2, 0, -0.30001780793026E-03),
				ijn(2, 1, 0.47661393906987E-04),
				ijn(2, 3, -0.44141845330846E-05),
				ijn(2, 17, -0.72694996297594E-15),
				ijn(3, -4, -0.31679644845054E-04),
				ijn(3, 0, -0.28270797985312E-05),
				ijn(3, 6, -0.85205128120103E-09),
				ijn(4, -5, -0.22425281908000E-05),
				ijn(4, -2, -0.65171222895601E-06),
				ijn(4, 10, -0.14341729937924E-12),
				ijn(5, -8, -0.40516996860117E-06),
				ijn(8, -11, -0.12734301741641E-08),
				ijn(8, -6, -0.17424871230634E-09),
				ijn(21, -29, -0.68762131295531E-18),
				ijn(23, -31, 0.14478307828521E-19),
				ijn(29, -38, 0.26335781662795E-22),
				ijn(30, -39, -0.11947622640071E-22),
				ijn(31, -40, 0.18228094581404E-23),
				ijn(32, -41, -0.93537087292458E-25)	]
	// Region2
	pt0_r2 = [	jn(0, -0.96927686500217E+01),
				jn(1, 0.10086655968018E+02),
				jn(-5, -0.56087911283020E-02),
				jn(-4, 0.71452738081455E-01),
				jn(-3, -0.40710498223928E+00),
				jn(-2, 0.14240819171444E+01),
				jn(-1, -0.43839511319450E+01),
				jn(2, -0.28408632460772E+00),
				jn(3, 0.21268463753307E-01)]
	pt1_r2 = [	ijn(1, 0, -0.17731742473213E-02),
				ijn(1, 1, -0.17834862292358E-01),
				ijn(1, 2, -0.45996013696365E-01),
				ijn(1, 3, -0.57581259083432E-01),
				ijn(1, 6, -0.50325278727930E-01),
				ijn(2, 1, -0.33032641670203E-04),
				ijn(2, 2, -0.18948987516315E-03),
				ijn(2, 4, -0.39392777243355E-02),
				ijn(2, 7, -0.43797295650573E-01),
				ijn(2, 36, -0.26674547914087E-04),
				ijn(3, 0, 0.20481737692309E-07),
				ijn(3, 1, 0.43870667284435E-06),
				ijn(3, 3, -0.32277677238570E-04),
				ijn(3, 6, -0.15033924542148E-02),
				ijn(3, 35, -0.40668253562649E-01),
				ijn(4, 1, -0.78847309559367E-09),
				ijn(4, 2, 0.12790717852285E-07),
				ijn(4, 3, 0.48225372718507E-06),
				ijn(5, 7, 0.22922076337661E-05),
				ijn(6, 3, -0.16714766451061E-10),
				ijn(6, 16, -0.21171472321355E-02),
				ijn(6, 35, -0.23895741934104E+02),
				ijn(7, 0, -0.59059564324270E-17),
				ijn(7, 11, -0.12621808899101E-05),
				ijn(7, 25, -0.38946842435739E-01),
				ijn(8, 8, 0.11256211360459E-10),
				ijn(8, 36, -0.82311340897998E+01),
				ijn(9, 13, 0.19809712802088E-07),
				ijn(10, 4, 0.10406965210174E-18),
				ijn(10, 10, -0.10234747095929E-12),
				ijn(10, 14, -0.10018179379511E-08),
				ijn(16, 29, -0.80882908646985E-10),
				ijn(16, 50, 0.10693031879409E+00),
				ijn(18, 57, -0.33662250574171E+00),
				ijn(20, 20, 0.89185845355421E-24),
				ijn(20, 35, 0.30629316876232E-12),
				ijn(20, 48, -0.42002467698208E-05),
				ijn(21, 21, -0.59056029685639E-25),
				ijn(22, 53, 0.37826947613457E-05),
				ijn(23, 39, -0.12768608934681E-14),
				ijn(24, 26, 0.73087610595061E-28),
				ijn(24, 40, 0.55414715350778E-16),
				ijn(24, 58, -0.94369707241210E-06)	]
	// Region3
	n1_r3 = 0.10658070028513E+01
	rt_r3 = [	ijn(0, 0, -0.15732845290239E+02),
				ijn(0, 1, 0.20944396974307E+02),
				ijn(0, 2, -0.76867707878716E+01),
				ijn(0, 7, 0.26185947787954E+01),
				ijn(0, 10, -0.28080781148620E+01),
				ijn(0, 12, 0.12053369696517E+01),
				ijn(0, 23, -0.84566812812502E-02),
				ijn(1, 2, -0.12654315477714E+01),
				ijn(1, 6, -0.11524407806681E+01),
				ijn(1, 15, 0.88521043984318E+00),
				ijn(1, 17, -0.64207765181607E+00),
				ijn(2, 0, 0.38493460186671E+00),
				ijn(2, 2, -0.85214708824206E+00),
				ijn(2, 6, 0.48972281541877E+01),
				ijn(2, 7, -0.30502617256965E+01),
				ijn(2, 22, 0.39420536879154E-01),
				ijn(2, 26, 0.12558408424308E+00),
				ijn(3, 0, -0.27999329698710E+00),
				ijn(3, 2, 0.13899799569460E+01),
				ijn(3, 4, -0.20189915023570E+01),
				ijn(3, 16, -0.82147637173963E-02),
				ijn(3, 26, -0.47596035734923E+00),
				ijn(4, 0, 0.43984074473500E-01),
				ijn(4, 2, -0.44476435428739E+00),
				ijn(4, 4, 0.90572070719733E+00),
				ijn(4, 26, 0.70522450087967E+00),
				ijn(5, 1, 0.10770512626332E+00),
				ijn(5, 3, -0.32913623258954E+00),
				ijn(5, 26, -0.50871062041158E+00),
				ijn(6, 0, -0.22175400873096E-01),
				ijn(6, 2, 0.94260751665092E-01),
				ijn(6, 26, 0.16436278447961E+00),
				ijn(7, 2, -0.13503372241348E-01),
				ijn(8, 26, -0.14834345352472E-01),
				ijn(9, 2, 0.57922953628084E-03),
				ijn(9, 26, 0.32308904703711E-02),
				ijn(10, 0, 0.80964802996215E-04),
				ijn(10, 1, -0.16557679795037E-03),
				ijn(11, 26, -0.44923899061815E-04)]
	// Region4 :
	pt_r4 = [	0.11670521452767E+04, 
				-0.72421316703206E+06,
				-0.17073846940092E+02,
				0.12020824702470E+05,
				-0.32325550322333E+07,
				0.14915108613530E+02,
				-0.48232657361591E+04,
				0.40511340542057E+06,
				-0.23855557567849E+00,
				-0.65017534844798E+03 ]
	// Region4 : rhof(T), rhog(T)
	t1_r4 = [1.99274064, 1.09965342, -0.510839303, -1.75493479, -45.5170352, -6.74694450E+05]
	t2_r4 = [-2.03150240, -2.68302940, -5.38626492, -17.2991605, -44.7586581, -63.9201063]
	// Region5
	pt_r5 = [	// Ideal Part
				ijn(0, 0, -1.3179983674201e1),
				ijn(0, 1, 6.8540841634434),
				ijn(0, -3, -2.4805148933466E-2),
				ijn(0, -2, 3.6901534980333E-1),
				ijn(0, -1, -3.1161318213925),
				ijn(0, 2, -3.2961626538917E-1),
				// Residual Part
				ijn(1, 1, 0.15736404855259E-2),
				ijn(1, 2, 0.90153761673944E-3),
				ijn(1, 3, -0.50270077677648E-2),
				ijn(2, 3, 0.22440037409485E-5),
				ijn(2, 9, -0.41163275453471E-5),
				ijn(3, 7, 0.37919454822955E-7)]
)

//****************************************************************
// CONST FOR `BOUNDS` EQUATIONS
//****************************************************************
const (
	//  Region 1 3 boundary h(s) calculation
	s_b13 = [	ijn(0, 0, 0.913965547600543), 
				ijn(1, -2, -0.430944856041991E-4), 
				ijn(1, 2, 0.603235694765419e2),
				ijn(3, -12, 0.117518273082168E-17), 
				ijn(5, -4, 0.220000904781292),
				ijn(6, -3, -0.690815545851641e2)]

	//  Region 1 4 boundary h(s) calculation
	s_b14 = [	ijn(0, 0, 0.913965547600543), 
				ijn(1, -2, -0.430944856041991E-4), 
				ijn(1, 2, 0.603235694765419e2),
				ijn(3, -12, 0.117518273082168E-17), 
				ijn(5, -4, 0.220000904781292),
				ijn(6, -3, -0.690815545851641e2)]
	// Region 2 : subregions
	hp_b2bc = [9.0584278514723e2, -6.7955786399241E-1, 1.2809002730136E-4,
				2.6526571908428e3, 4.5257578905948]	
    hs_b2ab = [-0.349898083432139e4, 0.257560716905876e4, -0.421073558227969e3, 0.276349063799944e2]
	//  Region 2 3 boundary p(T), T(p) calculation
	tp_b23 = [	0.34805185628969E+03, -0.11671859879975E+01, 0.10192970039326E-02, 
				0.57254459862746E+03, 0.13918839778870E+02]
	hs_b23 = [	ijn(-12, 10, 6.29096260829810E-04),
				ijn(-10, 8, -8.23453502583165E-04),
				ijn(-8, 3, 5.15446951519474E-08),
				ijn(-4, 4, -1.17565945784945E+00),
				ijn(-3, 3, 3.48519684726192E+00),
				ijn(-2, -6, -5.07837382408313E-12),
				ijn(-2, 2, -2.84637670005479E+00),
				ijn(-2, 3, -2.36092263939673E+00),
				ijn(-2, 4, 6.01492324973779E+00),
				ijn(0, 0, 1.48039650824546E+00),
				ijn(1, -3, 3.60075182221907E-04),
				ijn(1, -2, -1.26700045009952E-02),
				ijn(1, 10, -1.22184332521413E+06),
				ijn(3, -2, 1.49276502463272E-01),
				ijn(3, -1, 6.98733471798484E-01),
				ijn(5, -5, -2.52207040114321E-02),
				ijn(6, -6, 1.47151930985213E-02),
				ijn(6, -3, -1.08618917681849E+00),
				ijn(8, -8, -9.36875039816322E-04),
				ijn(8, -2, 8.19877897570217E+01),
				ijn(8, -1, -1.82041861521835E+02),
				ijn(12, -12, 2.61907376402688E-06),
				ijn(12, -1, -2.91626417025961E+04),
				ijn(14, -12, 1.40660774926165E-05),
				ijn(14, 1, 7.83237062349385E+06)]
	// Region 3 (Saturated Line) : b3_psat_h, 
	h_b3 = [	ijn(0, 0, 6.00073641753024E-01), 
				ijn(1, 1, -9.36203654849857E+00), 
				ijn(1, 3, 2.46590798594147E+01), 
				ijn(1, 4, -1.07014222858224E+02), 
				ijn(1, 36, -9.15821315805768E+13), 
				ijn(5, 3, -8.62332011700662E+03), 
				ijn(7, 0, -2.35837344740032E+01), 
				ijn(8, 24, 2.52304969384128E+17), 
				ijn(14, 16, -3.89718771997719E+18), 
				ijn(20, 16, -3.33775713645296E+22), 
				ijn(22, 3, 3.56499469636328E+10), 
				ijn(24, 18, -1.48547544720641E+26), 
				ijn(28, 8, 3.30611514838798E+18), 
				ijn(36, 24, 8.13641294467829E+37)]		
	// Region 3 (Saturated Line) : b3_psat_s, 
	s_b3 = [	ijn(1 , 1 , -1.29727445396014E+01), 
				ijn(1 , 32 , -2.24595125848403E+15), 
				ijn(4 , 7 , 1.77466741801846E+06), 
				ijn(12 , 4 , 7.17079349571538E+09), 
				ijn(12 , 14 , -3.78829107169011E+17), 
				ijn(16 , 36 , -9.55586736431328E+34), 
				ijn(24 , 10 , 1.87269814676188E+23), 
				ijn(28 , 0 , 1.19254746466473E+11), 
				ijn(32 , 18 , 1.10649277244882E+36)]
)
